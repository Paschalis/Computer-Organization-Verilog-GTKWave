module submodule_hw_8_c_or(
    output wire F1,
    input wire A,B
);
or U0 (F1, A, B);
endmodule    