module submodule_hw_8_c_not(
    output wire F1,
    input wire A
);
not U0 (F1, A);
endmodule
