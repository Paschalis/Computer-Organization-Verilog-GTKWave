`timescale 1ns / 1ps

module demultiplexer(
    in,
    s0,s1,s2,
    d0,d1,d2,d3,d4,d5,d6,d7);
input in,s0,s1,s2;
output d0,d1,d2,d3,d4,d5,d6,d7;
assign  d0=(in & ~s2 & ~s1 &~s0),
        d1=(in & ~s2 & ~s1 &s0),
        d2=(in & ~s2 & s1 &~s0),
        d3=(in & ~s2 & s1 &s0),
        d4=(in & s2 & ~s1 &~s0),
        d5=(in & s2 & ~s1 &s0),
        d6=(in & s2 & s1 &~s0),
        d7=(in & s2 & s1 &s0);
endmodule