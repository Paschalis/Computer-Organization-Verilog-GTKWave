module submodule_hw_8_b_or(
    output wire F1,
    input wire A, B, C, D, E, F, G, H 
);    
or U0 (F1, A, B, C, D, E, F, G, H);
endmodule