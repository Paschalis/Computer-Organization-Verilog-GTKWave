module submodule_hw_8_a(
    output wire y,
    input wire a,b,c,d
);

nand U0 (y, a, b, c, d);
endmodule

