module submodule_hw_8_b_and(
    output wire F1,
    input wire A, B, C, D 
);    
and U0 (F1, A, B, C, D);
endmodule