module submodule_xor(
    output wire XOR,
    input wire A,B
);
xor U0 (XOR, A, B);
endmodule