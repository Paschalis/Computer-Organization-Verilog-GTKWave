module submodule_hw_8_c_xor(
    output wire F1,
    input wire A,B
);
xor U0 (F1, A, B);
endmodule
